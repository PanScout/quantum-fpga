library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
--use work.fixed.ALL;
--use IEEE.fixed_pkg.ALL;
use work.fixed_pkg.ALL;

use work.qTypes.all;

entity Ceiling_Of_Log2 is
    port (
        scalar : in cfixedHigh;
        result : out cfixedHigh
    );
end Ceiling_Of_Log2;

architecture Structural of Ceiling_Of_Log2 is
    -- Threshold constants for 2^(n-1) where n is output value
constant TH_25 : fixedHigh := "0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
constant TH_24 : fixedHigh := "0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
constant TH_23 : fixedHigh := "0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
constant TH_22 : fixedHigh := "0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
constant TH_21 : fixedHigh := "0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
constant TH_20 : fixedHigh := "0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
constant TH_19 : fixedHigh := "0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
constant TH_18 : fixedHigh := "0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
constant TH_17 : fixedHigh := "0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000";
constant TH_16 : fixedHigh := "0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
constant TH_15 : fixedHigh := "0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000";
constant TH_14 : fixedHigh := "0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
constant TH_13 : fixedHigh := "0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000";
constant TH_12 : fixedHigh := "0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000";
constant TH_11 : fixedHigh := "0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000";
constant TH_10 : fixedHigh := "0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
constant TH_9 : fixedHigh := "0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
constant TH_8 : fixedHigh := "0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000";
constant TH_7 : fixedHigh := "0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000";
constant TH_6 : fixedHigh := "0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000";
constant TH_5 : fixedHigh := "0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000";
constant TH_4 : fixedHigh := "0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
constant TH_3 : fixedHigh := "0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
constant TH_2 : fixedHigh := "0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
constant TH_1 : fixedHigh := "0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
begin
    -- Ceiling log2 calculation using priority-encoded thresholds
    result.re <= 
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001" when scalar.re >= TH_25 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000" when scalar.re >= TH_24 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111" when scalar.re >= TH_23 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110" when scalar.re >= TH_22 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101" when scalar.re >= TH_21 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100" when scalar.re >= TH_20 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011" when scalar.re >= TH_19 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010" when scalar.re >= TH_18 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001" when scalar.re >= TH_17 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000" when scalar.re >= TH_16 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111" when scalar.re >= TH_15 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110" when scalar.re >= TH_14 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101" when scalar.re >= TH_13 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100" when scalar.re >= TH_12 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011" when scalar.re >= TH_11 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010" when scalar.re >= TH_10 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001" when scalar.re >= TH_9 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000" when scalar.re >= TH_8 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111" when scalar.re >= TH_7 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110" when scalar.re >= TH_6 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101" when scalar.re >= TH_5 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100" when scalar.re >= TH_4 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011" when scalar.re >= TH_3 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010" when scalar.re >= TH_2 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001" when scalar.re >= TH_1 else
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

    -- Imaginary component always zero
    result.im <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
end Structural;
