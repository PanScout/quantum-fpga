library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
--use work.fixed64.ALL;
--use IEEE.fixed_pkg.ALL;
use work.fixed_pkg.ALL;

use work.qTypes.all;

entity Ceiling_Of_Log2 is
    port (
        scalar : in cfixed64;
        result : out cfixed64
    );
end Ceiling_Of_Log2;

architecture Structural of Ceiling_Of_Log2 is
    -- Threshold constants for 2^(n-1) where n is output value
--constant TH_25 : fixed64 := "0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_24 : fixed64 := "0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_23 : fixed64 := "0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_22 : fixed64 := "0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_21 : fixed64 := "0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_20 : fixed64 := "0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_19 : fixed64 := "0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_18 : fixed64 := "0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_17 : fixed64 := "0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_16 : fixed64 := "0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_15 : fixed64 := "0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_14 : fixed64 := "0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_13 : fixed64 := "0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_12 : fixed64 := "0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_11 : fixed64 := "0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_10 : fixed64 := "0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_9 : fixed64 := "0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_8 : fixed64 := "0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_7 : fixed64 := "0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_6 : fixed64 := "0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_5 : fixed64 := "0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_4 : fixed64 := "0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_3 : fixed64 := "0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_2 : fixed64 := "0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
--constant TH_1 : fixed64 := "0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
--constant TH_0 : fixed64 := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";	      

     constant TH_25 : fixed64 := to_sfixed(2**24, fixed64'high, fixed64'low);
     constant TH_24 : fixed64 := to_sfixed(2**23, fixed64'high, fixed64'low);
     constant TH_23 : fixed64 := to_sfixed(2**22, fixed64'high, fixed64'low);
     constant TH_22 : fixed64 := to_sfixed(2**21, fixed64'high, fixed64'low);
     constant TH_21 : fixed64 := to_sfixed(2**20, fixed64'high, fixed64'low);
     constant TH_20 : fixed64 := to_sfixed(2**19, fixed64'high, fixed64'low);
     constant TH_19 : fixed64 := to_sfixed(2**18, fixed64'high, fixed64'low);
     constant TH_18 : fixed64 := to_sfixed(2**17, fixed64'high, fixed64'low);
     constant TH_17 : fixed64 := to_sfixed(2**16, fixed64'high, fixed64'low);
     constant TH_16 : fixed64 := to_sfixed(2**15, fixed64'high, fixed64'low);
     constant TH_15 : fixed64 := to_sfixed(2**14, fixed64'high, fixed64'low);
     constant TH_14 : fixed64 := to_sfixed(2**13, fixed64'high, fixed64'low);
     constant TH_13 : fixed64 := to_sfixed(2**12, fixed64'high, fixed64'low);
     constant TH_12 : fixed64 := to_sfixed(2**11, fixed64'high, fixed64'low);
     constant TH_11 : fixed64 := to_sfixed(2**10, fixed64'high, fixed64'low);
     constant TH_10 : fixed64 := to_sfixed(2**9,  fixed64'high, fixed64'low);
     constant TH_9  : fixed64 := to_sfixed(2**8,  fixed64'high, fixed64'low);
     constant TH_8  : fixed64 := to_sfixed(2**7,  fixed64'high, fixed64'low);
     constant TH_7  : fixed64 := to_sfixed(2**6,  fixed64'high, fixed64'low);
     constant TH_6  : fixed64 := to_sfixed(2**5,  fixed64'high, fixed64'low);
     constant TH_5  : fixed64 := to_sfixed(2**4,  fixed64'high, fixed64'low);
     constant TH_4  : fixed64 := to_sfixed(2**3,  fixed64'high, fixed64'low);
     constant TH_3  : fixed64 := to_sfixed(2**2,  fixed64'high, fixed64'low);
     constant TH_2  : fixed64 := to_sfixed(2**1,  fixed64'high, fixed64'low);
     constant TH_1  : fixed64 := to_sfixed(2**0,  fixed64'high, fixed64'low);

begin
    -- Ceiling log2 calculation using priority-encoded thresholds
    result.re <= 
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001" when scalar.re >= TH_25 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000" when scalar.re >= TH_24 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111" when scalar.re >= TH_23 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110" when scalar.re >= TH_22 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101" when scalar.re >= TH_21 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100" when scalar.re >= TH_20 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011" when scalar.re >= TH_19 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010" when scalar.re >= TH_18 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001" when scalar.re >= TH_17 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000" when scalar.re >= TH_16 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111" when scalar.re >= TH_15 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110" when scalar.re >= TH_14 else
----"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101" when scalar.re >= TH_13 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100" when scalar.re >= TH_12 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011" when scalar.re >= TH_11 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010" when scalar.re >= TH_10 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001" when scalar.re >= TH_9 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000" when scalar.re >= TH_8 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111" when scalar.re >= TH_7 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110" when scalar.re >= TH_6 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101" when scalar.re >= TH_5 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100" when scalar.re >= TH_4 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011" when scalar.re >= TH_3 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010" when scalar.re >= TH_2 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001" when scalar.re >= TH_1 else
--"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

         to_sfixed(25, fixed64'high, fixed64'low) when scalar.re >= TH_25 else
         to_sfixed(24, fixed64'high, fixed64'low) when scalar.re >= TH_24 else
         to_sfixed(23, fixed64'high, fixed64'low) when scalar.re >= TH_23 else
         to_sfixed(22, fixed64'high, fixed64'low) when scalar.re >= TH_22 else
         to_sfixed(21, fixed64'high, fixed64'low) when scalar.re >= TH_21 else
         to_sfixed(20, fixed64'high, fixed64'low) when scalar.re >= TH_20 else
         to_sfixed(19, fixed64'high, fixed64'low) when scalar.re >= TH_19 else
         to_sfixed(18, fixed64'high, fixed64'low) when scalar.re >= TH_18 else
         to_sfixed(17, fixed64'high, fixed64'low) when scalar.re >= TH_17 else
         to_sfixed(16, fixed64'high, fixed64'low) when scalar.re >= TH_16 else
         to_sfixed(15, fixed64'high, fixed64'low) when scalar.re >= TH_15 else
         to_sfixed(14, fixed64'high, fixed64'low) when scalar.re >= TH_14 else
         to_sfixed(13, fixed64'high, fixed64'low) when scalar.re >= TH_13 else
         to_sfixed(12, fixed64'high, fixed64'low) when scalar.re >= TH_12 else
         to_sfixed(11, fixed64'high, fixed64'low) when scalar.re >= TH_11 else
         to_sfixed(10, fixed64'high, fixed64'low) when scalar.re >= TH_10 else
         to_sfixed(9,  fixed64'high, fixed64'low) when scalar.re >= TH_9  else
         to_sfixed(8,  fixed64'high, fixed64'low) when scalar.re >= TH_8  else
         to_sfixed(7,  fixed64'high, fixed64'low) when scalar.re >= TH_7  else
         to_sfixed(6,  fixed64'high, fixed64'low) when scalar.re >= TH_6  else
         to_sfixed(5,  fixed64'high, fixed64'low) when scalar.re >= TH_5  else
         to_sfixed(4,  fixed64'high, fixed64'low) when scalar.re >= TH_4  else
         to_sfixed(3,  fixed64'high, fixed64'low) when scalar.re >= TH_3  else
         to_sfixed(2,  fixed64'high, fixed64'low) when scalar.re >= TH_2  else
         to_sfixed(1,  fixed64'high, fixed64'low) when scalar.re >= TH_1  else
         to_sfixed(0,  fixed64'high, fixed64'low);
    -- Imaginary component always zero
    result.im <= "0000000000000000000000000000000000000000000000000000000000000000";
    --result.im <= to_sfixed(0.0, fixed64'high, fixed64'low);
end Structural;
