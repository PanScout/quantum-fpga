library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.fixed_pkg.ALL;
use work.qTypes.ALL;

entity Pade_Denominator is
    Port (
        B : in  cmatrixHigh;
        P : out cmatrixHigh
    );
end Pade_Denominator;

architecture Structural of Pade_Denominator is

    ----------------------------------------------------------------------------
    -- Component Declarations
    ----------------------------------------------------------------------------
    component Matrix_Plus_Scalar_High is
        port (
            input_cMatrixH : in  cmatrixHigh;
            scalar         : in  cfixedHigh;
            output_cMatrixH: out cmatrixHigh
        );
    end component;
    
    component Matrix_By_Matrix_Multiplication_High is
        port (
            A : in  cmatrixHigh;
            B : in  cmatrixHigh;
            C : out cmatrixHigh
        );
    end component;
    
    ----------------------------------------------------------------------------
    -- Constant Coefficient Declarations for Numerator (all imaginary parts are zero)
    ----------------------------------------------------------------------------
    constant coeff1 : cfixedHigh := ( re => "1111111111111111111111111111111111111111111101001100000000000000000000000000000000000000000000000000000000000000000",
                                      im => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
    constant coeff2 : cfixedHigh := ( re => "0000000000000000000000000000000000000001111011110000000000000000000000000000000000000000000000000000000000000000000",
                                      im => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
    constant coeff3 : cfixedHigh := ( re => "1111111111111111111111111111111111001001110111000000000000000000000000000000000000000000000000000000000000000000000",
                                      im => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
    constant coeff4 : cfixedHigh := ( re => "0000000000000000000000000000010000011111101111100000000000000000000000000000000000000000000000000000000000000000000",
				      im => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
    constant coeff5 : cfixedHigh := ( re => "1111111111111111111111111100011001000011100111000000000000000000000000000000000000000000000000000000000000000000000",
                                      im => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
    constant coeff6 : cfixedHigh := ( re => "0000000000000000000000100100000101011011111010000000000000000000000000000000000000000000000000000000000000000000000",
                                      im => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
    constant coeff7 : cfixedHigh := ( re => "1111111111111111111100001000100011110111100000000000000000000000000000000000000000000000000000000000000000000000000",
                                      im => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
    constant coeff8 : cfixedHigh := ( re => "0000000000000000010000011011100111100100001000000000000000000000000000000000000000000000000000000000000000000000000",
                                      im => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
    constant coeff9 : cfixedHigh := ( re => "1111111111111111011111001000110000110111110000000000000000000000000000000000000000000000000000000000000000000000000",
                                      im => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
                                      

    ----------------------------------------------------------------------------
    -- Signal Declarations for Intermediate Results
    ----------------------------------------------------------------------------
    signal T0, T1, T2, T3, T4, T5, T6, T7, T8 : cmatrixHigh;
    signal M1, M2, M3, M4, M5, M6, M7, M8       : cmatrixHigh;

begin

    -- T0 = B + coeff1  (i.e. B + 90)
    U0: Matrix_Plus_Scalar_High
        port map (
            input_cMatrixH => B,
            scalar         => coeff1,
            output_cMatrixH=> T0
        );
    
    -- M1 = T0 * B
    U1: Matrix_By_Matrix_Multiplication_High
        port map (
            A => T0,
            B => B,
            C => M1
        );
    
    -- T1 = M1 + coeff2
    U2: Matrix_Plus_Scalar_High
        port map (
            input_cMatrixH => M1,
            scalar         => coeff2,
            output_cMatrixH=> T1
        );
    
    -- M2 = T1 * B
    U3: Matrix_By_Matrix_Multiplication_High
        port map (
            A => T1,
            B => B,
            C => M2
        );
    
    -- T2 = M2 + coeff3
    U4: Matrix_Plus_Scalar_High
        port map (
            input_cMatrixH => M2,
            scalar         => coeff3,
            output_cMatrixH=> T2
        );
    
    -- M3 = T2 * B
    U5: Matrix_By_Matrix_Multiplication_High
        port map (
            A => T2,
            B => B,
            C => M3
        );
    
    -- T3 = M3 + coeff4
    U6: Matrix_Plus_Scalar_High
        port map (
            input_cMatrixH => M3,
            scalar         => coeff4,
            output_cMatrixH=> T3
        );
    
    -- M4 = T3 * B
    U7: Matrix_By_Matrix_Multiplication_High
        port map (
            A => T3,
            B => B,
            C => M4
        );
    
    -- T4 = M4 + coeff5
    U8: Matrix_Plus_Scalar_High
        port map (
            input_cMatrixH => M4,
            scalar         => coeff5,
            output_cMatrixH=> T4
        );
    
    -- M5 = T4 * B
    U9: Matrix_By_Matrix_Multiplication_High
        port map (
            A => T4,
            B => B,
            C => M5
        );
    
    -- T5 = M5 + coeff6
    U10: Matrix_Plus_Scalar_High
        port map (
            input_cMatrixH => M5,
            scalar         => coeff6,
            output_cMatrixH=> T5
        );
    
    -- M6 = T5 * B
    U11: Matrix_By_Matrix_Multiplication_High
        port map (
            A => T5,
            B => B,
            C => M6
        );
    
    -- T6 = M6 + coeff7
    U12: Matrix_Plus_Scalar_High
        port map (
            input_cMatrixH => M6,
            scalar         => coeff7,
            output_cMatrixH=> T6
        );
    
    -- M7 = T6 * B
    U13: Matrix_By_Matrix_Multiplication_High
        port map (
            A => T6,
            B => B,
            C => M7
        );
    
    -- T7 = M7 + coeff8
    U14: Matrix_Plus_Scalar_High
        port map (
            input_cMatrixH => M7,
            scalar         => coeff8,
            output_cMatrixH=> T7
        );
    
    -- M8 = T7 * B
    U15: Matrix_By_Matrix_Multiplication_High
        port map (
            A => T7,
            B => B,
            C => M8
        );
    
    -- T8 = M8 + coeff9  --> Final result
    U16: Matrix_Plus_Scalar_High
        port map (
            input_cMatrixH => M8,
            scalar         => coeff9,
            output_cMatrixH=> T8
        );

   P <= T8;

end Structural;
